-----------------------------------------------------------
--This file is automatically generated for the network given as
--X = [15,5,7,12,16,20,27,2,6,7,10,11,14,17,18,20,25,2,3,15,26,15,18,24,26,1,10,11,14,15,16,23,25,26,4,5,6,11,12,19,1,3,4,5,6,12,14,18,19,20,24,26,2,4,5,10,11,12,14,18,19,27,4,14,18,27,5,10,12,13,19,20,24,26,4,10,18,7,8,10,22,25,26,1,2,4,11,15,2,7,12,20,21,25,27,1,8,17,22,4,6,8,9,10,15,25,1,4,15,24,25,1,5,6,10,14,15,16,17,27,9,12,13,18,27,2,4,5,6,10,14,25,1,2,3,6,10,11,15,21,24,25,27,1,5,8,15,18,20,22,27,4,4,5,9,12,24,2,3,7,10,12,14,21,4,7,17,18,21,24,28,29,30]
--Xn= [1,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,4,4,4,4,5,5,5,5,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,10,10,10,10,11,11,11,11,11,11,11,11,12,12,12,13,13,13,13,13,13,14,14,14,14,14,15,15,15,15,15,15,15,16,16,16,16,17,17,17,17,17,17,17,18,18,18,18,18,19,19,19,19,19,19,19,19,19,20,20,20,20,20,21,21,21,21,21,21,21,22,22,22,22,22,22,22,22,22,22,22,23,23,23,23,23,23,23,23,24,25,25,25,25,25,26,26,26,26,26,26,26,27,27,27,27,27,27,1,2,3]
--Tau=[1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1]
--W=[3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,3.00000,6.00000,3.00000,6.00000,3.00000,3.00000,3.00000,6.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,6.00000,3.00000,6.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,-5.00000,-2.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-2.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,6.00000,3.00000,3.00000,3.00000,3.00000,6.00000,3.00000,6.00000,3.00000,6.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,6.00000,3.00000,3.00000,3.00000,6.00000,3.00000,6.00000,3.00000,3.00000,6.00000,6.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,6.00000,3.00000,3.00000,3.00000,3.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-2.00000,-5.00000,-5.00000,-5.00000,-5.00000,-2.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-2.00000,-5.00000,-5.00000,-5.00000,-2.00000,-5.00000,3.00000,3.00000,3.00000,6.00000,3.00000,3.00000,-5.00000,-2.00000,-5.00000,-5.00000,-5.00000,-5.00000,-2.00000,3.00000,3.00000,3.00000,3.00000,6.00000,3.00000,1.00000,1.00000,1.00000]
--inputNeurons=[1,2,3]
--inputWeights=[1.00000,1.00000,1.00000]
--inputDelays=[1,1,1]
--outputNeurons=[1,2,3,4,5,6,7,8,9,10]
-----------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

library ieee_proposed;
use ieee_proposed.fixed_pkg.all;
use ieee_proposed.math_utility_pkg.all;

library work;
use work.myTypes.all;
use work.all;


entity Network is
port (clk,globalRst : in std_logic;
        spikeIn: in std_logic_vector(3 downto 1);
        spikeOut: out std_logic_vector(10 downto 1));
end entity;

architecture arch of Network is
component neuron is
        -- neuron parameters
        generic( Nsyn : natural :=3;
           D : integerArray:=(2,3,4);
           W : realArray:=(0.5, 0.2, 0.3);
           alpha_w :real :=1.0;
           beta_w  :real :=0.1;
           alpha_v1:real :=0.98;
           alpha_v2:real :=0.9333;
           alpha_V :real :=0.98;
           alpha_A :real :=0.98;
           beta_1  :real :=0.286;
           beta_2  :real :=1.0;
           beta_A  :real :=-0.1;
           V_th :real :=1.0);

       port ( inputSpikes : in std_logic_vector(Nsyn downto 1):=(others=>'0');
              outputSpike : out std_logic:='0';
              globalRst,clk : in std_logic:='0';
              Iapp : in fp:=to_sfixed(0,fp_int,fp_frac));
end component;


   --Define common neuron parameters
   constant alpha_w  :real :=1.00000;
   constant alpha_v1 :real :=0.98000;
   constant alpha_v2 :real :=0.93330;
   constant alpha_V  :real :=0.98000;
   constant alpha_A  :real :=0.98000;
   constant beta_1   :real :=0.28600;
   constant beta_2   :real :=1.00000;
   constant beta_A   :real :=0.10000;
   constant beta_w   :real :=0.10000;
   constant V_th     :real :=1.00000;


   --Define interconnection delays for each neuron 
   constant D1 :integerArray :=(1,1);
   constant D2 :integerArray :=(1,1,1,1,1,1,1);
   constant D3 :integerArray :=(1,1,1,1,1,1,1,1,1,1,1);
   constant D4 :integerArray :=(1,1,1,1);
   constant D5 :integerArray :=(1,1,1,1);
   constant D6 :integerArray :=(1,1,1,1,1,1,1,1,1);
   constant D7 :integerArray :=(1,1,1,1,1,1);
   constant D8 :integerArray :=(1,1,1,1,1,1,1,1,1,1,1,1);
   constant D9 :integerArray :=(1,1,1,1,1,1,1,1,1,1);
   constant D10 :integerArray :=(1,1,1,1);
   constant D11 :integerArray :=(1,1,1,1,1,1,1,1);
   constant D12 :integerArray :=(1,1,1);
   constant D13 :integerArray :=(1,1,1,1,1,1);
   constant D14 :integerArray :=(1,1,1,1,1);
   constant D15 :integerArray :=(1,1,1,1,1,1,1);
   constant D16 :integerArray :=(1,1,1,1);
   constant D17 :integerArray :=(1,1,1,1,1,1,1);
   constant D18 :integerArray :=(1,1,1,1,1);
   constant D19 :integerArray :=(1,1,1,1,1,1,1,1,1);
   constant D20 :integerArray :=(1,1,1,1,1);
   constant D21 :integerArray :=(1,1,1,1,1,1,1);
   constant D22 :integerArray :=(1,1,1,1,1,1,1,1,1,1,1);
   constant D23 :integerArray :=(1,1,1,1,1,1,1,1);
   constant D24 :integerArray :=(1,1);
   constant D25 :integerArray :=(1,1,1,1,1);
   constant D26 :integerArray :=(1,1,1,1,1,1,1);
   constant D27 :integerArray :=(1,1,1,1,1,1);


   --Define initial Weights for each neuron
   constant W1 :realArray :=(3.00000,1.00000);
   constant W2 :realArray :=(3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,1.00000);
   constant W3 :realArray :=(-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,1.00000);
   constant W4 :realArray :=(3.00000,6.00000,3.00000,6.00000);
   constant W5 :realArray :=(3.00000,3.00000,3.00000,6.00000);
   constant W6 :realArray :=(3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,6.00000,3.00000,6.00000);
   constant W7 :realArray :=(3.00000,3.00000,3.00000,3.00000,3.00000,3.00000);
   constant W8 :realArray :=(-5.00000,-2.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-2.00000);
   constant W9 :realArray :=(-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000);
   constant W10 :realArray :=(3.00000,3.00000,3.00000,3.00000);
   constant W11 :realArray :=(3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,6.00000);
   constant W12 :realArray :=(3.00000,3.00000,3.00000);
   constant W13 :realArray :=(3.00000,6.00000,3.00000,6.00000,3.00000,6.00000);
   constant W14 :realArray :=(3.00000,3.00000,3.00000,3.00000,3.00000);
   constant W15 :realArray :=(3.00000,3.00000,3.00000,3.00000,6.00000,3.00000,3.00000);
   constant W16 :realArray :=(3.00000,6.00000,3.00000,6.00000);
   constant W17 :realArray :=(3.00000,3.00000,6.00000,6.00000,3.00000,3.00000,3.00000);
   constant W18 :realArray :=(3.00000,3.00000,3.00000,3.00000,3.00000);
   constant W19 :realArray :=(3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000,3.00000);
   constant W20 :realArray :=(6.00000,3.00000,3.00000,3.00000,3.00000);
   constant W21 :realArray :=(-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000,-5.00000);
   constant W22 :realArray :=(-5.00000,-5.00000,-2.00000,-5.00000,-5.00000,-5.00000,-5.00000,-2.00000,-5.00000,-5.00000,-5.00000);
   constant W23 :realArray :=(-5.00000,-5.00000,-2.00000,-5.00000,-5.00000,-5.00000,-2.00000,-5.00000);
   constant W24 :realArray :=(3.00000,1.0);
   constant W25 :realArray :=(3.00000,3.00000,6.00000,3.00000,3.00000);
   constant W26 :realArray :=(-5.00000,-2.00000,-5.00000,-5.00000,-5.00000,-5.00000,-2.00000);
   constant W27 :realArray :=(3.00000,3.00000,3.00000,3.00000,6.00000,3.00000);


   --Define interconnection signals
   signal synapseSpike1: std_logic_vector(2 downto 1):=(others=>'0');
   signal synapseSpike2: std_logic_vector(7 downto 1):=(others=>'0');
   signal synapseSpike3: std_logic_vector(11 downto 1):=(others=>'0');
   signal synapseSpike4: std_logic_vector(4 downto 1):=(others=>'0');
   signal synapseSpike5: std_logic_vector(4 downto 1):=(others=>'0');
   signal synapseSpike6: std_logic_vector(9 downto 1):=(others=>'0');
   signal synapseSpike7: std_logic_vector(6 downto 1):=(others=>'0');
   signal synapseSpike8: std_logic_vector(12 downto 1):=(others=>'0');
   signal synapseSpike9: std_logic_vector(10 downto 1):=(others=>'0');
   signal synapseSpike10: std_logic_vector(4 downto 1):=(others=>'0');
   signal synapseSpike11: std_logic_vector(8 downto 1):=(others=>'0');
   signal synapseSpike12: std_logic_vector(3 downto 1):=(others=>'0');
   signal synapseSpike13: std_logic_vector(6 downto 1):=(others=>'0');
   signal synapseSpike14: std_logic_vector(5 downto 1):=(others=>'0');
   signal synapseSpike15: std_logic_vector(7 downto 1):=(others=>'0');
   signal synapseSpike16: std_logic_vector(4 downto 1):=(others=>'0');
   signal synapseSpike17: std_logic_vector(7 downto 1):=(others=>'0');
   signal synapseSpike18: std_logic_vector(5 downto 1):=(others=>'0');
   signal synapseSpike19: std_logic_vector(9 downto 1):=(others=>'0');
   signal synapseSpike20: std_logic_vector(5 downto 1):=(others=>'0');
   signal synapseSpike21: std_logic_vector(7 downto 1):=(others=>'0');
   signal synapseSpike22: std_logic_vector(11 downto 1):=(others=>'0');
   signal synapseSpike23: std_logic_vector(8 downto 1):=(others=>'0');
   signal synapseSpike24: std_logic_vector(1 downto 1):=(others=>'0');
   signal synapseSpike25: std_logic_vector(5 downto 1):=(others=>'0');
   signal synapseSpike26: std_logic_vector(7 downto 1):=(others=>'0');
   signal synapseSpike27: std_logic_vector(6 downto 1):=(others=>'0');

   signal Iapp : fp_array(27 downto 1):=(others=>to_sfixed(0.0,fp_int,fp_frac));
   signal neuronSpike: std_logic_vector(30 downto 1):=(others=>'0');
begin


   --Generate Neurons
	N1 :  neuron generic map(Nsyn=>2,D=>D1,W=>W1,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(1),inputSpikes=>synapseSpike1,outputSpike=>neuronSpike(1),globalRst=>globalRst,clk=>clk);
	N2 :  neuron generic map(Nsyn=>7,D=>D2,W=>W2,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(2),inputSpikes=>synapseSpike2,outputSpike=>neuronSpike(2),globalRst=>globalRst,clk=>clk);
	N3 :  neuron generic map(Nsyn=>11,D=>D3,W=>W3,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(3),inputSpikes=>synapseSpike3,outputSpike=>neuronSpike(3),globalRst=>globalRst,clk=>clk);
	N4 :  neuron generic map(Nsyn=>4,D=>D4,W=>W4,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(4),inputSpikes=>synapseSpike4,outputSpike=>neuronSpike(4),globalRst=>globalRst,clk=>clk);
	N5 :  neuron generic map(Nsyn=>4,D=>D5,W=>W5,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(5),inputSpikes=>synapseSpike5,outputSpike=>neuronSpike(5),globalRst=>globalRst,clk=>clk);
	N6 :  neuron generic map(Nsyn=>9,D=>D6,W=>W6,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(6),inputSpikes=>synapseSpike6,outputSpike=>neuronSpike(6),globalRst=>globalRst,clk=>clk);
	N7 :  neuron generic map(Nsyn=>6,D=>D7,W=>W7,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(7),inputSpikes=>synapseSpike7,outputSpike=>neuronSpike(7),globalRst=>globalRst,clk=>clk);
	N8 :  neuron generic map(Nsyn=>12,D=>D8,W=>W8,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(8),inputSpikes=>synapseSpike8,outputSpike=>neuronSpike(8),globalRst=>globalRst,clk=>clk);
	N9 :  neuron generic map(Nsyn=>10,D=>D9,W=>W9,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(9),inputSpikes=>synapseSpike9,outputSpike=>neuronSpike(9),globalRst=>globalRst,clk=>clk);
	N10 :  neuron generic map(Nsyn=>4,D=>D10,W=>W10,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(10),inputSpikes=>synapseSpike10,outputSpike=>neuronSpike(10),globalRst=>globalRst,clk=>clk);
	N11 :  neuron generic map(Nsyn=>8,D=>D11,W=>W11,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(11),inputSpikes=>synapseSpike11,outputSpike=>neuronSpike(11),globalRst=>globalRst,clk=>clk);
	N12 :  neuron generic map(Nsyn=>3,D=>D12,W=>W12,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(12),inputSpikes=>synapseSpike12,outputSpike=>neuronSpike(12),globalRst=>globalRst,clk=>clk);
	N13 :  neuron generic map(Nsyn=>6,D=>D13,W=>W13,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(13),inputSpikes=>synapseSpike13,outputSpike=>neuronSpike(13),globalRst=>globalRst,clk=>clk);
	N14 :  neuron generic map(Nsyn=>5,D=>D14,W=>W14,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(14),inputSpikes=>synapseSpike14,outputSpike=>neuronSpike(14),globalRst=>globalRst,clk=>clk);
	N15 :  neuron generic map(Nsyn=>7,D=>D15,W=>W15,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(15),inputSpikes=>synapseSpike15,outputSpike=>neuronSpike(15),globalRst=>globalRst,clk=>clk);
	N16 :  neuron generic map(Nsyn=>4,D=>D16,W=>W16,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(16),inputSpikes=>synapseSpike16,outputSpike=>neuronSpike(16),globalRst=>globalRst,clk=>clk);
	N17 :  neuron generic map(Nsyn=>7,D=>D17,W=>W17,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(17),inputSpikes=>synapseSpike17,outputSpike=>neuronSpike(17),globalRst=>globalRst,clk=>clk);
	N18 :  neuron generic map(Nsyn=>5,D=>D18,W=>W18,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(18),inputSpikes=>synapseSpike18,outputSpike=>neuronSpike(18),globalRst=>globalRst,clk=>clk);
	N19 :  neuron generic map(Nsyn=>9,D=>D19,W=>W19,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(19),inputSpikes=>synapseSpike19,outputSpike=>neuronSpike(19),globalRst=>globalRst,clk=>clk);
	N20 :  neuron generic map(Nsyn=>5,D=>D20,W=>W20,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(20),inputSpikes=>synapseSpike20,outputSpike=>neuronSpike(20),globalRst=>globalRst,clk=>clk);
	N21 :  neuron generic map(Nsyn=>7,D=>D21,W=>W21,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(21),inputSpikes=>synapseSpike21,outputSpike=>neuronSpike(21),globalRst=>globalRst,clk=>clk);
	N22 :  neuron generic map(Nsyn=>11,D=>D22,W=>W22,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(22),inputSpikes=>synapseSpike22,outputSpike=>neuronSpike(22),globalRst=>globalRst,clk=>clk);
	N23 :  neuron generic map(Nsyn=>8,D=>D23,W=>W23,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(23),inputSpikes=>synapseSpike23,outputSpike=>neuronSpike(23),globalRst=>globalRst,clk=>clk);
	N24 :  neuron generic map(Nsyn=>1,D=>D24,W=>W24,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(24),inputSpikes=>synapseSpike24,outputSpike=>neuronSpike(24),globalRst=>globalRst,clk=>clk);
	N25 :  neuron generic map(Nsyn=>5,D=>D25,W=>W25,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(25),inputSpikes=>synapseSpike25,outputSpike=>neuronSpike(25),globalRst=>globalRst,clk=>clk);
	N26 :  neuron generic map(Nsyn=>7,D=>D26,W=>W26,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(26),inputSpikes=>synapseSpike26,outputSpike=>neuronSpike(26),globalRst=>globalRst,clk=>clk);
	N27 :  neuron generic map(Nsyn=>6,D=>D27,W=>W27,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(27),inputSpikes=>synapseSpike27,outputSpike=>neuronSpike(27),globalRst=>globalRst,clk=>clk);


   --Map Synapses
   synapseSpike1(1)<=neuronSpike(15);
   synapseSpike1(2)<=neuronSpike(28);
   synapseSpike2(1)<=neuronSpike(5);
   synapseSpike2(2)<=neuronSpike(7);
   synapseSpike2(3)<=neuronSpike(12);
   synapseSpike2(4)<=neuronSpike(16);
   synapseSpike2(5)<=neuronSpike(20);
   synapseSpike2(6)<=neuronSpike(27);
   synapseSpike2(7)<=neuronSpike(29);
   synapseSpike3(1)<=neuronSpike(2);
   synapseSpike3(2)<=neuronSpike(6);
   synapseSpike3(3)<=neuronSpike(7);
   synapseSpike3(4)<=neuronSpike(10);
   synapseSpike3(5)<=neuronSpike(11);
   synapseSpike3(6)<=neuronSpike(14);
   synapseSpike3(7)<=neuronSpike(17);
   synapseSpike3(8)<=neuronSpike(18);
   synapseSpike3(9)<=neuronSpike(20);
   synapseSpike3(10)<=neuronSpike(25);
   synapseSpike3(11)<=neuronSpike(30);
   synapseSpike4(1)<=neuronSpike(2);
   synapseSpike4(2)<=neuronSpike(3);
   synapseSpike4(3)<=neuronSpike(15);
   synapseSpike4(4)<=neuronSpike(26);
   synapseSpike5(1)<=neuronSpike(15);
   synapseSpike5(2)<=neuronSpike(18);
   synapseSpike5(3)<=neuronSpike(24);
   synapseSpike5(4)<=neuronSpike(26);
   synapseSpike6(1)<=neuronSpike(1);
   synapseSpike6(2)<=neuronSpike(10);
   synapseSpike6(3)<=neuronSpike(11);
   synapseSpike6(4)<=neuronSpike(14);
   synapseSpike6(5)<=neuronSpike(15);
   synapseSpike6(6)<=neuronSpike(16);
   synapseSpike6(7)<=neuronSpike(23);
   synapseSpike6(8)<=neuronSpike(25);
   synapseSpike6(9)<=neuronSpike(26);
   synapseSpike7(1)<=neuronSpike(4);
   synapseSpike7(2)<=neuronSpike(5);
   synapseSpike7(3)<=neuronSpike(6);
   synapseSpike7(4)<=neuronSpike(11);
   synapseSpike7(5)<=neuronSpike(12);
   synapseSpike7(6)<=neuronSpike(19);
   synapseSpike8(1)<=neuronSpike(1);
   synapseSpike8(2)<=neuronSpike(3);
   synapseSpike8(3)<=neuronSpike(4);
   synapseSpike8(4)<=neuronSpike(5);
   synapseSpike8(5)<=neuronSpike(6);
   synapseSpike8(6)<=neuronSpike(12);
   synapseSpike8(7)<=neuronSpike(14);
   synapseSpike8(8)<=neuronSpike(18);
   synapseSpike8(9)<=neuronSpike(19);
   synapseSpike8(10)<=neuronSpike(20);
   synapseSpike8(11)<=neuronSpike(24);
   synapseSpike8(12)<=neuronSpike(26);
   synapseSpike9(1)<=neuronSpike(2);
   synapseSpike9(2)<=neuronSpike(4);
   synapseSpike9(3)<=neuronSpike(5);
   synapseSpike9(4)<=neuronSpike(10);
   synapseSpike9(5)<=neuronSpike(11);
   synapseSpike9(6)<=neuronSpike(12);
   synapseSpike9(7)<=neuronSpike(14);
   synapseSpike9(8)<=neuronSpike(18);
   synapseSpike9(9)<=neuronSpike(19);
   synapseSpike9(10)<=neuronSpike(27);
   synapseSpike10(1)<=neuronSpike(4);
   synapseSpike10(2)<=neuronSpike(14);
   synapseSpike10(3)<=neuronSpike(18);
   synapseSpike10(4)<=neuronSpike(27);
   synapseSpike11(1)<=neuronSpike(5);
   synapseSpike11(2)<=neuronSpike(10);
   synapseSpike11(3)<=neuronSpike(12);
   synapseSpike11(4)<=neuronSpike(13);
   synapseSpike11(5)<=neuronSpike(19);
   synapseSpike11(6)<=neuronSpike(20);
   synapseSpike11(7)<=neuronSpike(24);
   synapseSpike11(8)<=neuronSpike(26);
   synapseSpike12(1)<=neuronSpike(4);
   synapseSpike12(2)<=neuronSpike(10);
   synapseSpike12(3)<=neuronSpike(18);
   synapseSpike13(1)<=neuronSpike(7);
   synapseSpike13(2)<=neuronSpike(8);
   synapseSpike13(3)<=neuronSpike(10);
   synapseSpike13(4)<=neuronSpike(22);
   synapseSpike13(5)<=neuronSpike(25);
   synapseSpike13(6)<=neuronSpike(26);
   synapseSpike14(1)<=neuronSpike(1);
   synapseSpike14(2)<=neuronSpike(2);
   synapseSpike14(3)<=neuronSpike(4);
   synapseSpike14(4)<=neuronSpike(11);
   synapseSpike14(5)<=neuronSpike(15);
   synapseSpike15(1)<=neuronSpike(2);
   synapseSpike15(2)<=neuronSpike(7);
   synapseSpike15(3)<=neuronSpike(12);
   synapseSpike15(4)<=neuronSpike(20);
   synapseSpike15(5)<=neuronSpike(21);
   synapseSpike15(6)<=neuronSpike(25);
   synapseSpike15(7)<=neuronSpike(27);
   synapseSpike16(1)<=neuronSpike(1);
   synapseSpike16(2)<=neuronSpike(8);
   synapseSpike16(3)<=neuronSpike(17);
   synapseSpike16(4)<=neuronSpike(22);
   synapseSpike17(1)<=neuronSpike(4);
   synapseSpike17(2)<=neuronSpike(6);
   synapseSpike17(3)<=neuronSpike(8);
   synapseSpike17(4)<=neuronSpike(9);
   synapseSpike17(5)<=neuronSpike(10);
   synapseSpike17(6)<=neuronSpike(15);
   synapseSpike17(7)<=neuronSpike(25);
   synapseSpike18(1)<=neuronSpike(1);
   synapseSpike18(2)<=neuronSpike(4);
   synapseSpike18(3)<=neuronSpike(15);
   synapseSpike18(4)<=neuronSpike(24);
   synapseSpike18(5)<=neuronSpike(25);
   synapseSpike19(1)<=neuronSpike(1);
   synapseSpike19(2)<=neuronSpike(5);
   synapseSpike19(3)<=neuronSpike(6);
   synapseSpike19(4)<=neuronSpike(10);
   synapseSpike19(5)<=neuronSpike(14);
   synapseSpike19(6)<=neuronSpike(15);
   synapseSpike19(7)<=neuronSpike(16);
   synapseSpike19(8)<=neuronSpike(17);
   synapseSpike19(9)<=neuronSpike(27);
   synapseSpike20(1)<=neuronSpike(9);
   synapseSpike20(2)<=neuronSpike(12);
   synapseSpike20(3)<=neuronSpike(13);
   synapseSpike20(4)<=neuronSpike(18);
   synapseSpike20(5)<=neuronSpike(27);
   synapseSpike21(1)<=neuronSpike(2);
   synapseSpike21(2)<=neuronSpike(4);
   synapseSpike21(3)<=neuronSpike(5);
   synapseSpike21(4)<=neuronSpike(6);
   synapseSpike21(5)<=neuronSpike(10);
   synapseSpike21(6)<=neuronSpike(14);
   synapseSpike21(7)<=neuronSpike(25);
   synapseSpike22(1)<=neuronSpike(1);
   synapseSpike22(2)<=neuronSpike(2);
   synapseSpike22(3)<=neuronSpike(3);
   synapseSpike22(4)<=neuronSpike(6);
   synapseSpike22(5)<=neuronSpike(10);
   synapseSpike22(6)<=neuronSpike(11);
   synapseSpike22(7)<=neuronSpike(15);
   synapseSpike22(8)<=neuronSpike(21);
   synapseSpike22(9)<=neuronSpike(24);
   synapseSpike22(10)<=neuronSpike(25);
   synapseSpike22(11)<=neuronSpike(27);
   synapseSpike23(1)<=neuronSpike(1);
   synapseSpike23(2)<=neuronSpike(5);
   synapseSpike23(3)<=neuronSpike(8);
   synapseSpike23(4)<=neuronSpike(15);
   synapseSpike23(5)<=neuronSpike(18);
   synapseSpike23(6)<=neuronSpike(20);
   synapseSpike23(7)<=neuronSpike(22);
   synapseSpike23(8)<=neuronSpike(27);
   synapseSpike24(1)<=neuronSpike(4);
   synapseSpike25(1)<=neuronSpike(4);
   synapseSpike25(2)<=neuronSpike(5);
   synapseSpike25(3)<=neuronSpike(9);
   synapseSpike25(4)<=neuronSpike(12);
   synapseSpike25(5)<=neuronSpike(24);
   synapseSpike26(1)<=neuronSpike(2);
   synapseSpike26(2)<=neuronSpike(3);
   synapseSpike26(3)<=neuronSpike(7);
   synapseSpike26(4)<=neuronSpike(10);
   synapseSpike26(5)<=neuronSpike(12);
   synapseSpike26(6)<=neuronSpike(14);
   synapseSpike26(7)<=neuronSpike(21);
   synapseSpike27(1)<=neuronSpike(4);
   synapseSpike27(2)<=neuronSpike(7);
   synapseSpike27(3)<=neuronSpike(17);
   synapseSpike27(4)<=neuronSpike(18);
   synapseSpike27(5)<=neuronSpike(21);
   synapseSpike27(6)<=neuronSpike(24);


   --Map Inputs from external world 
   neuronSpike(28)<=spikeIn(1);
   neuronSpike(29)<=spikeIn(2);
   neuronSpike(30)<=spikeIn(3);


   --Map Outputs to external world 
   spikeOut(1)<=neuronSpike(1);
   spikeOut(2)<=neuronSpike(2);
   spikeOut(3)<=neuronSpike(3);
   spikeOut(4)<=neuronSpike(4);
   spikeOut(5)<=neuronSpike(5);
   spikeOut(6)<=neuronSpike(6);
   spikeOut(7)<=neuronSpike(7);
   spikeOut(8)<=neuronSpike(8);
   spikeOut(9)<=neuronSpike(9);
   spikeOut(10)<=neuronSpike(10);
end arch;
