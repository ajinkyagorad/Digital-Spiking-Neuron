-----------------------------------------------------------
--This file is automatically generated for the network given as
--X = [1,1,1,2,2,2,3,3,3,5,6,7]
--Xn= [2,3,4,1,3,4,1,2,4,1,2,3]
--Tau=[1,2,3,4,5,6,7,8,9,1,1,1]
--W=[0.10000,0.20000,0.30000,0.40000,0.50000,0.60000,0.70000,0.80000,0.90000,1.00000,1.00000,1.00000]
--inputNeurons=[1,2,3]
--inputWeights=[1.00000,1.00000,1.00000]
--inputDelays=[1,1,1]
--outputNeurons=[4]
-----------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

library ieee_proposed;
use ieee_proposed.fixed_pkg.all;
use ieee_proposed.math_utility_pkg.all;

library work;
use work.myTypes.all;
use work.all;


entity Network is
port (clk,globalRst : in std_logic;
        spikeIn: in std_logic_vector(3 downto 1);
        spikeOut: out std_logic_vector(1 downto 1));
end entity;

architecture arch of Network is
component neuron is
        -- neuron parameters
        generic( Nsyn : natural :=3;
           D : integerArray:=(2,3,4);
           W : realArray:=(0.5, 0.2, 0.3);
           alpha_w :real :=1.0;
           beta_w  :real :=0.1;
           alpha_v1:real :=0.98;
           alpha_v2:real :=0.9333;
           alpha_V :real :=0.98;
           alpha_A :real :=0.98;
           beta_1  :real :=0.286;
           beta_2  :real :=1.0;
           beta_A  :real :=-0.1;
           V_th :real :=1.0);

       port ( inputSpikes : in std_logic_vector(Nsyn downto 1):=(others=>'0');
              outputSpike : out std_logic:='0';
              globalRst,clk : in std_logic:='0';
              Iapp : in fp:=to_sfixed(0,fp_int,fp_frac));
end component;


   --Define common neuron parameters
   constant alpha_w  :real :=1.00000;
   constant alpha_v1 :real :=0.98000;
   constant alpha_v2 :real :=0.93330;
   constant alpha_V  :real :=0.98000;
   constant alpha_A  :real :=0.98000;
   constant beta_1   :real :=0.28600;
   constant beta_2   :real :=1.00000;
   constant beta_A   :real :=0.10000;
   constant beta_w   :real :=0.10000;
   constant V_th     :real :=1.00000;


   --Define interconnection delays for each neuron 
   constant D1 :integerArray :=(4,7,1);
   constant D2 :integerArray :=(1,8,1);
   constant D3 :integerArray :=(2,5,1);
   constant D4 :integerArray :=(3,6,9);


   --Define initial Weights for each neuron
   constant W1 :realArray :=(0.40000,0.70000,1.00000);
   constant W2 :realArray :=(0.10000,0.80000,1.00000);
   constant W3 :realArray :=(0.20000,0.50000,1.00000);
   constant W4 :realArray :=(0.30000,0.60000,0.90000);


   --Define interconnection signals
   signal synapseSpike1: std_logic_vector(3 downto 1):=(others=>'0');
   signal synapseSpike2: std_logic_vector(3 downto 1):=(others=>'0');
   signal synapseSpike3: std_logic_vector(3 downto 1):=(others=>'0');
   signal synapseSpike4: std_logic_vector(3 downto 1):=(others=>'0');

   signal Iapp : fp_array(4 downto 1):=(others=>to_sfixed(0.0,fp_int,fp_frac));
   signal neuronSpike: std_logic_vector(7 downto 1):=(others=>'0');
begin


   --Generate Neurons
	N1 :  neuron generic map(Nsyn=>3,D=>D1,W=>W1,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(1),inputSpikes=>synapseSpike1,outputSpike=>neuronSpike(1),globalRst=>globalRst,clk=>clk);
	N2 :  neuron generic map(Nsyn=>3,D=>D2,W=>W2,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(2),inputSpikes=>synapseSpike2,outputSpike=>neuronSpike(2),globalRst=>globalRst,clk=>clk);
	N3 :  neuron generic map(Nsyn=>3,D=>D3,W=>W3,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(3),inputSpikes=>synapseSpike3,outputSpike=>neuronSpike(3),globalRst=>globalRst,clk=>clk);
	N4 :  neuron generic map(Nsyn=>3,D=>D4,W=>W4,alpha_V=>alpha_V,alpha_v1=>alpha_v1,alpha_v2=>alpha_v2,alpha_A=>alpha_A,alpha_w=>alpha_w,beta_1=>beta_1,beta_2=>beta_2,beta_A=>beta_A,beta_w=>beta_w)
           port map(Iapp=>Iapp(4),inputSpikes=>synapseSpike4,outputSpike=>neuronSpike(4),globalRst=>globalRst,clk=>clk);


   --Map Synapses
   synapseSpike1(1)<=neuronSpike(2);
   synapseSpike1(2)<=neuronSpike(3);
   synapseSpike1(3)<=neuronSpike(5);
   synapseSpike2(1)<=neuronSpike(1);
   synapseSpike2(2)<=neuronSpike(3);
   synapseSpike2(3)<=neuronSpike(6);
   synapseSpike3(1)<=neuronSpike(1);
   synapseSpike3(2)<=neuronSpike(2);
   synapseSpike3(3)<=neuronSpike(7);
   synapseSpike4(1)<=neuronSpike(1);
   synapseSpike4(2)<=neuronSpike(2);
   synapseSpike4(3)<=neuronSpike(3);


   --Map Inputs from external world 
   neuronSpike(5)<=spikeIn(1);
   neuronSpike(6)<=spikeIn(2);
   neuronSpike(7)<=spikeIn(3);


   --Map Outputs to external world 
   spikeOut(1)<=neuronSpike(4);
end arch;
